module decoder(IR, NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD,
					SUB, INAC, CLAC, AND, OR, XOR, NOT);

	input [7:0] IR;

	output reg NOP;
	output reg LDAC;
	output reg STAC;
	output reg MVAC;
	output reg MOVR;
	output reg JUMP;
	output reg JMPZ;
	output reg JPNZ;
	output reg ADD;
	output reg SUB;
	output reg INAC;
	output reg CLAC;
	output reg AND;
	output reg OR;
	output reg XOR;
	output reg NOT;
	
	always @(*)
	begin
		if ( ~(IR[7]|IR[6]|IR[5]|IR[4]) == 0)
				{NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_0000_0000_0000;
		else
			begin
				case(IR[3:0])
					4'b0000: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b1000_0000_0000_0000;
					4'b0001: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0100_0000_0000_0000;
					4'b0010: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0010_0000_0000_0000;
					4'b0011: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0001_0000_0000_0000;
					4'b0100: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_1000_0000_0000;
					4'b0101: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_0100_0000_0000;
					4'b0110: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_0010_0000_0000;
					4'b0111: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_0001_0000_0000;
					4'b1000: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_0000_1000_0000;
					4'b1001: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_0000_0100_0000;
					4'b1010: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_0000_0010_0000;
					4'b1011: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_0000_0001_0000;
					4'b1100: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_0000_0000_1000;
					4'b1101: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_0000_0000_0100;
					4'b1110: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_0000_0000_0010;
					4'b1111: {NOP, LDAC, STAC, MVAC, MOVR, JUMP, JMPZ, JPNZ, ADD, SUB, INAC, CLAC, AND, OR, XOR, NOT} = 16'b0000_0000_0000_0001;
				endcase
			end
	end
	
endmodule
				